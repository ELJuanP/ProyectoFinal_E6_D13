`timescale 1ns/1ns
module And(
	input A,
	input B,
	output C
);

assign C = A & B;
endmodule