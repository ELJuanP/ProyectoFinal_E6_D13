`timescale 1ns/1ns
module Adder1 (
	input [3:0]A,
	output[3:0]B
);

assign B = A + 4;
endmodule
