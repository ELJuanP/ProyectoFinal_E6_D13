'timescale 1ns/1ns

module Alu-Control;
	input [5:0]OpCode;
	output MemToReg;
	output MemToWrite;
	output ALUOp;
	output RegToWrite;

wire c1, c3;
reg c2, c4;

assign c3 = ALUOp
 endmodule
